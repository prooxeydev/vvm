module releases

pub struct Assets {
pub:
	id int
	name string
}