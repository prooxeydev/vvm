module releases

struct Release {
pub:
	id int
	name string
	assets []Assets
}